library ieee;
use ieee.std_logic_1164.all;

ENTITY ProcessadorDidatico IS
	PORT(
		Clock , Reset : IN BIT
	);
END ProcessadorDidatico;

ARCHITECTURE ProcessadorDidatico_Arch OF ProcessadorDidatico IS
	BEGIN
END ProcessadorDidatico_Arch;